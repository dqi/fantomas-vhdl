library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;
use ieee.std_logic_unsigned.all;

entity fantomas_lbox is
	port (
		a1 : in std_logic_vector(7 downto 0);
		a2 : in std_logic_vector(7 downto 0);
		o : out std_logic_vector(15 downto 0)
	);
end entity fantomas_lbox;

architecture behav of fantomas_lbox is
  -----------------------------------------------------------------------------
  -- Type definitions
  -----------------------------------------------------------------------------
  subtype ByteInt is integer range 0 to 65335; type ByteArray is array (0 to 255) of ByteInt;
  -----------------------------------------------------------------------------
  -- Constants
  -----------------------------------------------------------------------------
  constant LBOX1 : ByteArray := (
  0, 49151, 28304, 53615, 16695, 65224, 12199, 36952, 54600, 27319, 48088, 1063,
  38015, 11136, 64239, 17680, 21142, 60777, 15366, 33785, 5025, 44126, 32049,
  49870, 34782, 14369, 59726, 22193, 50921, 30998, 43129, 6022, 53635, 28284,
  48915, 236, 37044, 12107, 65060, 16859, 1227, 47924, 27227, 54692, 17916,
  64003, 11116, 38035, 33557, 15594, 60805, 21114, 49698, 32221, 44210, 4941,
  22109, 59810, 14541, 34610, 5994, 43157, 31226, 50693, 49841, 32078, 44065,
  5086, 33670, 15481, 60694, 21225, 6137, 43014, 31081, 50838, 22222, 59697,
  14430, 34721, 36903, 12248, 65207, 16712, 53520, 28399, 49024, 127, 17775,
  64144, 11263, 37888, 1112, 48039, 27336, 54583, 4914, 44237, 32162, 49757,
  20997, 60922, 15509, 33642, 50810, 31109, 43242, 5909, 34637, 14514, 59869,
  22050, 16804, 65115, 12084, 37067, 147, 49004, 28163, 53756, 38124, 11027,
  64124, 17795, 54747, 27172, 47947, 1204, 18796, 63123, 10236, 38915, 2139,
  47012, 26315, 55604, 39972, 9179, 62132, 19787, 56595, 25324, 45955, 3196,
  7162, 41989, 30058, 51861, 23245, 58674, 13405, 35746, 52914, 29005, 40994,
  8157, 36741, 12410, 57621, 24298, 39151, 10000, 63103, 18816, 55768, 26151,
  46920, 2231, 19879, 62040, 9015, 40136, 3216, 45935, 25088, 56831, 51833,
  30086, 42217, 6934, 35662, 13489, 58846, 23073, 7985, 41166, 29089, 52830,
  24070, 57849, 12438, 36713, 35805, 13346, 58701, 23218, 51946, 29973, 42106,
  7045, 24213, 57706, 12293, 36858, 8098, 41053, 28978, 52941, 55627, 26292,
  47067, 2084, 39036, 10115, 63212, 18707, 3075, 46076, 25235, 56684, 19764,
  62155, 9124, 40027, 23134, 58785, 13518, 35633, 7017, 42134, 30201, 51718,
  36630, 12521, 57734, 24185, 52769, 29150, 41137, 8014, 2248, 46903, 26200,
  55719, 18943, 62976, 10095, 39056, 56704, 25215, 45840, 3311, 40119, 9032,
  61991, 19928
  );

  constant LBOX2 : ByteArray := (
  0, 29890, 54052, 42982, 52776, 47850, 7436, 27086, 26710, 7316, 47986, 53168,
  42622, 53948, 30042, 408, 58505, 36939, 14253, 17263, 10913, 24163, 63877,
  36167, 36063, 63517, 24571, 11065, 17143, 13877, 37331, 58641, 26681, 7419,
  47901, 53215, 42513, 53971, 30005, 503, 111, 29869, 54091, 42889, 52807,
  47749, 7523, 27041, 36016, 63602, 24468, 11094, 17048, 13914, 37308, 58750,
  58598, 36900, 14274, 17152, 10958, 24076, 63978, 36136, 24132, 10886, 36192,
  63906, 36972, 58542, 17224, 14218, 13842, 17104, 58678, 37364, 63546, 36088,
  11038, 24540, 47821, 52751, 27113, 7467, 29925, 39, 42945, 54019, 53915,
  42585, 447, 30077, 7347, 26737, 53143, 47957, 13949, 17087, 58713, 37275,
  63573, 35991, 11121, 24499, 24107, 10985, 36111, 63949, 36867, 58561, 17191,
  14309, 54004, 42550, 464, 29970, 7388, 26654, 53240, 47930, 47778, 52832,
  27014, 7492, 29834, 72, 42926, 54124, 24907, 5513, 45679, 50861, 44899, 56225,
  31815, 2181, 2333, 32223, 55865, 44795, 50997, 46071, 5137, 24787, 34242,
  61696, 22246, 8740, 19434, 16168, 39118, 60428, 60820, 39254, 16048, 19058,
  9148, 22398, 61592, 33882, 2418, 32176, 55894, 44692, 51034, 45976, 5246,
  24764, 24868, 5606, 45568, 50882, 44812, 56270, 31784, 2282, 60923, 39225,
  16095, 18973, 9171, 22289, 61687, 33845, 34221, 61807, 22153, 8779, 19333,
  16199, 39073, 60515, 16143, 19405, 60459, 39145, 61735, 34277, 8707, 22209,
  22361, 9115, 33917, 61631, 39281, 60851, 19029, 16023, 56198, 44868, 2210,
  31840, 5550, 24940, 50826, 45640, 46032, 50962, 24820, 5174, 32248, 2362,
  44764, 55838, 22326, 9204, 33810, 61648, 39198, 60892, 19002, 16120, 16224,
  19362, 60484, 39046, 61768, 34186, 8812, 22190, 46015, 51069, 24731, 5209,
  32151, 2389, 44723, 55921, 56297, 44843, 2253, 31759, 5569, 24835, 50917,
  45607
  );

begin
  process (a1, a2)
    variable r1 : std_logic_vector(15 downto 0);
    variable r2 : std_logic_vector(15 downto 0);
  begin
    r1 := std_logic_vector(to_unsigned(LBOX1(to_integer(unsigned(a1))), 16));
    r2 := std_logic_vector(to_unsigned(LBOX2(to_integer(unsigned(a2))), 16));
    o <= r1 xor r2;
  end process;
end architecture behav;
