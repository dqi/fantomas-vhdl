library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fantomas_transform is
  port (
    a : in std_logic_vector(127 downto 0);
    o : out std_logic_vector(127 downto 0)
  );
end entity fantomas_transform;

architecture behav of fantomas_transform is

  -- Variables
begin
  
end behav;
